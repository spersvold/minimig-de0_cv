// -*- mode: verilog; mode: font-lock; indent-tabs-mode: nil -*-
// vi: set et ts=3 sw=3 sts=3:
//
// Copyright 2006, 2007 Dennis van Weeren
//
// This file is part of Minimig
//
// Minimig is free software; you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation; either version 3 of the License, or
// (at your option) any later version.
//
// Minimig is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <http://www.gnu.org/licenses/>.
//
//
//
// This is the user IO module
//
//
// SP:
// 2016-03-24 - cleanup


module userio
  (
   input  wire        clk,                // bus clock
   input  wire        reset,              // reset
   input  wire        clk7_en,
   input  wire        clk7n_en,
   input  wire        c1,
   input  wire        c3,
   input  wire        sol,                // start of video line
   input  wire        sof,                // start of video frame
   input  wire        varbeamen,
   input  wire [ 8:1] reg_address_in,     // register adress inputs
   input  wire [15:0] data_in,            // bus data in
   output reg  [15:0] data_out,           // bus data out
   inout  wire        ps2mdat,            // mouse PS/2 data
   inout  wire        ps2mclk,            // mouse PS/2 clk
   output wire        _fire0,             // joystick 0 fire output (to CIA)
   output wire        _fire1,             // joystick 1 fire output (to CIA)
   input  wire        _fire0_dat,
   input  wire        _fire1_dat,
   input  wire        aflock,             // auto fire lock
   input  wire [ 7:0] _joy1,              // joystick 1 in (default mouse port)
   input  wire [ 7:0] _joy2,              // joystick 2 in (default joystick port)
   input  wire [ 5:0] mou_emu,
   input  wire [ 5:0] joy_emu,
   input  wire [ 7:0] osd_ctrl,           // OSD control (minimig->host, [menu,select,down,up])
   output wire        key_disable,        // disables Amiga keyboard while OSD is active
   input  wire        _scs,               // SPI enable
   input  wire        sdi,                // SPI data in
   output wire        sdo,                // SPI data out
   input  wire        sck,                // SPI clock
   output wire        osd_blank,          // osd overlay, normal video blank output
   output wire        osd_pixel,          // osd video pixel
   output wire [ 1:0] lr_filter,
   output wire [ 1:0] hr_filter,
   output wire [ 6:0] memory_config,
   output wire [ 4:0] chipset_config,
   output wire [ 3:0] floppy_config,
   output wire [ 1:0] scanline,
   output wire [ 1:0] dither,
   output wire [ 2:0] ide_config,
   output wire [ 3:0] cpu_config,
   output             usrrst,             // user reset from osd module
   output             cpurst,
   output             cpuhlt,
   output wire        fifo_full,
   // host
   output wire        host_cs,
   output wire [23:0] host_adr,
   output wire        host_we,
   output wire [ 1:0] host_bs,
   output wire [15:0] host_wdat,
   input  wire [15:0] host_rdat,
   input  wire        host_ack
   );

   // register names and adresses
   localparam JOY0DAT     = 9'h00a;
   localparam JOY1DAT     = 9'h00c;
   localparam SCRDAT      = 9'h1f0;
   localparam POTINP      = 9'h016;
   localparam POTGO       = 9'h034;
   localparam JOYTEST     = 9'h036;
   localparam KEY_MENU    = 8'h69;
   localparam KEY_ESC     = 8'h45;
   localparam KEY_ENTER   = 8'h44;
   localparam KEY_UP      = 8'h4C;
   localparam KEY_DOWN    = 8'h4D;
   localparam KEY_LEFT    = 8'h4F;
   localparam KEY_RIGHT   = 8'h4E;
   localparam KEY_PGUP    = 8'h6c;
   localparam KEY_PGDOWN  = 8'h6d;

   // local signals
   reg [ 7:0]         _sjoy1;           // synchronized joystick 1 signals
   reg [ 7:0]         _djoy1;           // synchronized joystick 1 signals
   reg [ 5:0]         _xjoy2;           // synchronized joystick 2 signals
   reg [ 7:0]         _tjoy2;           // synchronized joystick 2 signals
   reg [ 7:0]         _djoy2;           // synchronized joystick 2 signals
   wire [ 5:0]        _sjoy2;           // synchronized joystick 2 signals
   reg [15:0]         potreg;           // POTGO write
   wire [15:0]        mouse0dat;        // mouse counters
   wire [ 7:0]        mouse0scr;        // mouse scroller
   reg [15:0]         dmouse0dat;       // docking mouse counters
   reg [15:0]         dmouse1dat;       // docking mouse counters
   wire               _mleft;           // left mouse button
   wire               _mthird;          // middle mouse button
   wire               _mright;          // right mouse buttons
   reg                joy1enable;       // joystick 1 enable (mouse/joy switch)
   reg                joy2enable;       // joystick 2 enable when no osd
   wire               osd_enable;       // OSD display enable
   reg [ 7:0]         t_osd_ctrl;       // JB: osd control lines
   wire               test_load;        // load test value to mouse counter
   wire [15:0]        test_data;        // mouse counter test value
   wire [ 1:0]        autofire_config;
   reg [ 1:0]         autofire_cnt;
   wire               cd32pad;
   reg                autofire;
   reg                sel_autofire;     // select autofire and permanent fire
   reg [ 7:0]         cd32pad1_reg;
   reg [ 7:0]         cd32pad2_reg;

   //--------------------------------------------------------------------------------------
   //--------------------------------------------------------------------------------------

   // POTGO register
   always @ (posedge clk) begin
      if (clk7_en) begin
         if (reset)
           potreg <= #1 0;
         else if (reg_address_in[8:1]==POTGO[8:1])
           potreg[15:0] <= #1 data_in[15:0];
      end
   end

   // potcap reg
   reg  [4-1:0] potcap;
   always @ (posedge clk) begin
      if (clk7_en) begin
         if (reset)
           potcap <= #1 4'h0;
         else begin
            if (cd32pad && (potreg[15] && !potreg[14])) begin
               potcap[3] <= #1 cd32pad2_reg[7];
            end else begin
               if (!_sjoy2[5]) potcap[3] <= #1 1'b0;
               else if (potreg[15] & potreg[14]) potcap[3] <= #1 1'b1;
            end
            if (potreg[13]) potcap[2] <= #1 potreg[12];
            if (cd32pad && (potreg[11] && !potreg[10])) begin
               potcap[1] <= #1 cd32pad1_reg[7];
            end else begin
               if (!(_mright&_djoy1[5])) potcap[1] <= #1 1'b0;
               else if (potreg[11] & potreg[10]) potcap[1] <= #1 1'b1;
            end
            if (!_mthird) potcap[0] <= #1 1'b0;
            else if (potreg[ 9] & potreg[ 8]) potcap[0] <= #1 1'b1;
         end
      end
   end

   // cd32pad1 reg
   reg fire1_d;
   always @ (posedge clk) begin
      if (clk7_en) begin
         if (reset)
           fire1_d <= #1 1'b1;
         else
           fire1_d <= #1 _fire0_dat;
      end
   end
   wire cd32pad1_reg_load  = !(potreg[9] && !potreg[8]);
   wire cd32pad1_reg_shift = _fire0_dat && !fire1_d;
   always @ (posedge clk) begin
      if (clk7_en) begin
         if (reset)
           cd32pad1_reg <= #1 8'hff;
         else if (cd32pad1_reg_load)
           cd32pad1_reg <= #1 {_djoy1[5], _djoy1[4], _djoy1[6], _djoy1[7], 3'b111, 1'b1};
         else if (cd32pad1_reg_shift)
           cd32pad1_reg <= #1 {cd32pad1_reg[6:0], 1'b0};
      end
   end

   // cd32pad2 reg
   reg fire2_d;
   always @ (posedge clk) begin
      if (clk7_en) begin
         if (reset)
           fire2_d <= #1 1'b1;
         else
           fire2_d <= #1 _fire1_dat;
      end
   end
   wire cd32pad2_reg_load  = !(potreg[13] && !potreg[12]);
   wire cd32pad2_reg_shift = _fire1_dat && !fire2_d;
   always @ (posedge clk) begin
      if (clk7_en) begin
         if (reset)
           cd32pad2_reg <= #1 8'hff;
         else if (cd32pad2_reg_load)
           cd32pad2_reg <= #1 {_djoy2[5], _djoy2[4], _djoy2[6], _djoy2[7], 3'b111, 1'b1};
         else if (cd32pad2_reg_shift)
           cd32pad2_reg <= #1 {cd32pad2_reg[6:0], 1'b0};
      end
   end

   // autofire pulses generation
   always @ (posedge clk) begin
      if (clk7_en) begin
         if (sof)
           if (autofire_cnt == 1)
             autofire_cnt <= #1 autofire_config;
           else
             autofire_cnt <= #1 autofire_cnt - 2'd1;
      end
   end

   // autofire
   always @ (posedge clk) begin
      if (clk7_en) begin
         if (sof)
           if (autofire_config == 2'd0)
             autofire <= #1 1'b0;
           else if (autofire_cnt == 2'd1)
             autofire <= #1 ~autofire;
      end
   end

   // auto fire function toggle via capslock status
   always @ (posedge clk) begin
      if (clk7_en) begin
         sel_autofire <= #1 (~aflock ^ _xjoy2[4]) ? autofire : 1'b0;
      end
   end

   // input synchronization of external signals
   always @ (posedge clk) begin
      if (clk7_en) begin
         _sjoy1[7:0] <= #1 _joy1[7:0];
         _djoy1[7:0] <= #1 _sjoy1[7:0];
         _tjoy2[7:0] <= #1 _joy2[7:0] & {2'b11, joy_emu[5:0]};
         _djoy2[7:0] <= #1 _tjoy2[7:0];
         if (sof)
           _xjoy2[5:0] <= #1 _joy2[5:0] & joy_emu[5:0];
      end
   end

   // port 2 joystick disable in osd
   always @ (posedge clk) begin
      if (clk7_en) begin
         if (key_disable)
           joy2enable <= #1 0;
         else if (_xjoy2[5:0] == 6'b11_1111)
           joy2enable <= #1 1;
      end
   end

   // autofire is permanent active if enabled, can be overwritten any time by normal fire button
   assign _sjoy2[5:0] = joy2enable ? {_xjoy2[5], sel_autofire ^ _xjoy2[4], _xjoy2[3:0]} : 6'b11_1111;

   always @ (*) begin
      if (~joy2enable)
        if (~_xjoy2[5] || (~_xjoy2[3] && ~_xjoy2[2]))
          t_osd_ctrl = KEY_MENU;
        else if (~_xjoy2[4])
          t_osd_ctrl = KEY_ENTER;
        else if (~_xjoy2[3])
          t_osd_ctrl = KEY_UP;
        else if (~_xjoy2[2])
          t_osd_ctrl = KEY_DOWN;
        else if (~_xjoy2[1])
          t_osd_ctrl = KEY_LEFT;
        else if (~_xjoy2[0])
          t_osd_ctrl = KEY_RIGHT;
        else if (~_xjoy2[1] && ~_xjoy2[3])
          t_osd_ctrl = KEY_PGUP;
        else if (~_xjoy2[0] && ~_xjoy2[2])
          t_osd_ctrl = KEY_PGDOWN;
        else
          t_osd_ctrl = osd_ctrl;
      else
        t_osd_ctrl = osd_ctrl;
   end

   // port 1 automatic mouse/joystick switch
   always @ (posedge clk) begin
      if (clk7_en) begin
         if (!_mleft || reset)//when left mouse button pushed, switch to mouse (default)
           joy1enable = 0;
         else if (!_sjoy1[4])//when joystick 1 fire pushed, switch to joystick
           joy1enable = 1;
      end
   end

   // Port 1
   always @ (posedge clk) begin
      if (clk7_en) begin
         if (test_load)
           dmouse0dat[7:0] <= #1 8'h00;
         else if ((!_djoy1[0] && _sjoy1[0] && _sjoy1[2]) || (_djoy1[0] && !_sjoy1[0] && !_sjoy1[2]) || (!_djoy1[2] && _sjoy1[2] && !_sjoy1[0]) || (_djoy1[2] && !_sjoy1[2] && _sjoy1[0]))
           dmouse0dat[7:0] <= #1 dmouse0dat[7:0] + 1;
         else if ((!_djoy1[0] && _sjoy1[0] && !_sjoy1[2]) || (_djoy1[0] && !_sjoy1[0] && _sjoy1[2]) || (!_djoy1[2] && _sjoy1[2] && _sjoy1[0]) || (_djoy1[2] && !_sjoy1[2] && !_sjoy1[0]))
           dmouse0dat[7:0] <= #1 dmouse0dat[7:0] - 1;
         else
           dmouse0dat[1:0] <= #1 {!_djoy1[0], _djoy1[0] ^ _djoy1[2]};
      end
   end

   always @ (posedge clk) begin
      if (clk7_en) begin
         if (test_load)
           dmouse0dat[15:8] <= #1 8'h00;
         else if ((!_djoy1[1] && _sjoy1[1] && _sjoy1[3]) || (_djoy1[1] && !_sjoy1[1] && !_sjoy1[3]) || (!_djoy1[3] && _sjoy1[3] && !_sjoy1[1]) || (_djoy1[3] && !_sjoy1[3] && _sjoy1[1]))
           dmouse0dat[15:8] <= #1 dmouse0dat[15:8] + 1;
         else if ((!_djoy1[1] && _sjoy1[1] && !_sjoy1[3]) || (_djoy1[1] && !_sjoy1[1] && _sjoy1[3]) || (!_djoy1[3] && _sjoy1[3] && _sjoy1[1]) || (_djoy1[3] && !_sjoy1[3] && !_sjoy1[1]))
           dmouse0dat[15:8] <= #1 dmouse0dat[15:8] - 1;
         else
           dmouse0dat[9:8] <= #1 {!_djoy1[1], _djoy1[1] ^ _djoy1[3]};
      end
   end

   // Port 2
   always @ (posedge clk) begin
      if (clk7_en) begin
         if (test_load)
           dmouse1dat[7:2] <= #1 test_data[7:2];
         else if ((!_djoy2[0] && _tjoy2[0] && _tjoy2[2]) || (_djoy2[0] && !_tjoy2[0] && !_tjoy2[2]) || (!_djoy2[2] && _tjoy2[2] && !_tjoy2[0]) || (_djoy2[2] && !_tjoy2[2] && _tjoy2[0]))
           dmouse1dat[7:0] <= #1 dmouse1dat[7:0] + 1;
         else if ((!_djoy2[0] && _tjoy2[0] && !_tjoy2[2]) || (_djoy2[0] && !_tjoy2[0] && _tjoy2[2]) || (!_djoy2[2] && _tjoy2[2] && _tjoy2[0]) || (_djoy2[2] && !_tjoy2[2] && !_tjoy2[0]))
           dmouse1dat[7:0] <= #1 dmouse1dat[7:0] - 1;
         else
           dmouse1dat[1:0] <= #1 {!_djoy2[0], _djoy2[0] ^ _djoy2[2]};
      end
   end

   always @ (posedge clk) begin
      if (clk7_en) begin
         if (test_load)
           dmouse1dat[15:10] <= #1 test_data[15:10];
         else if ((!_djoy2[1] && _tjoy2[1] && _tjoy2[3]) || (_djoy2[1] && !_tjoy2[1] && !_tjoy2[3]) || (!_djoy2[3] && _tjoy2[3] && !_tjoy2[1]) || (_djoy2[3] && !_tjoy2[3] && _tjoy2[1]))
           dmouse1dat[15:8] <= #1 dmouse1dat[15:8] + 1;
         else if ((!_djoy2[1] && _tjoy2[1] && !_tjoy2[3]) || (_djoy2[1] && !_tjoy2[1] && _tjoy2[3]) || (!_djoy2[3] && _tjoy2[3] && _tjoy2[1]) || (_djoy2[3] && !_tjoy2[3] && !_tjoy2[1]))
           dmouse1dat[15:8] <= #1 dmouse1dat[15:8] - 1;
         else
           dmouse1dat[9:8] <= #1 {!_djoy2[1], _djoy2[1] ^ _djoy2[3]};
      end
   end

   //--------------------------------------------------------------------------------------
   //--------------------------------------------------------------------------------------

   // data output multiplexer
   always @(*) begin
      if ((reg_address_in[8:1]==JOY0DAT[8:1]) && joy1enable)//read port 1 joystick
        data_out[15:0] = {mouse0dat[15:10] + dmouse0dat[15:10],dmouse0dat[9:8],mouse0dat[7:2] + dmouse0dat[7:2],dmouse0dat[1:0]};
      else if (reg_address_in[8:1]==JOY0DAT[8:1])//read port 1 mouse
        data_out[15:0] = {mouse0dat[15:8] + dmouse0dat[15:8],mouse0dat[7:0] + dmouse0dat[7:0]};
      else if (reg_address_in[8:1]==JOY1DAT[8:1])//read port 2 joystick
        data_out[15:0] = dmouse1dat;
      else if (reg_address_in[8:1]==POTINP[8:1])//read mouse and joysticks extra buttons
        data_out[15:0] = {1'b0, potcap[3],
                          1'b0, potcap[2],
                          1'b0, potcap[1],
                          1'b0, potcap[0],
                          8'h00};
      else if (reg_address_in[8:1]==SCRDAT[8:1])//read mouse scroll wheel
        data_out[15:0] = {8'h00,mouse0scr};
      else
        data_out[15:0] = 16'h0000;
   end

   // assign fire outputs to cia A
   assign _fire0 = cd32pad && !cd32pad1_reg_load ? fire1_d : _sjoy1[4] & _mleft;
   assign _fire1 = cd32pad && !cd32pad2_reg_load ? fire2_d : _sjoy2[4];

   //JB: some trainers writes to JOYTEST register to reset current mouse counter
   assign test_load = reg_address_in[8:1]==JOYTEST[8:1] ? 1'b1 : 1'b0;
   assign test_data = data_in[15:0];

   //--------------------------------------------------------------------------------------
   //--------------------------------------------------------------------------------------

   //instantiate mouse controller
   userio_ps2mouse pm1
     (
      .clk        (clk),
      .clk7_en    (clk7_en),
      .reset      (reset),
      .ps2mdat    (ps2mdat),
      .ps2mclk    (ps2mclk),
      .mou_emu    (mou_emu),
      .sof        (sof),
      .zcount     (mouse0scr),
      .ycount     (mouse0dat[15:8]),
      .xcount     (mouse0dat[7:0]),
      ._mleft     (_mleft),
      ._mthird    (_mthird),
      ._mright    (_mright),
      .test_load  (test_load),
      .test_data  (test_data)
      );

   //--------------------------------------------------------------------------------------
   //--------------------------------------------------------------------------------------

   //instantiate osd controller
   userio_osd osd1
     (
      .clk              (clk),
      .clk7_en          (clk7_en),
      .clk7n_en         (clk7n_en),
      .reset            (reset),
      .c1               (c1),
      .c3               (c3),
      .sol              (sol),
      .sof              (sof),
      .varbeamen        (varbeamen),
      .osd_ctrl         (t_osd_ctrl),
      ._scs             (_scs),
      .sdi              (sdi),
      .sdo              (sdo),
      .sck              (sck),
      .osd_blank        (osd_blank),
      .osd_pixel        (osd_pixel),
      .osd_enable       (osd_enable),
      .key_disable      (key_disable),
      .lr_filter        (lr_filter),
      .hr_filter        (hr_filter),
      .memory_config    (memory_config),
      .chipset_config   (chipset_config),
      .floppy_config    (floppy_config),
      .scanline         (scanline),
      .dither           (dither),
      .ide_config       (ide_config),
      .cpu_config       (cpu_config),
      .autofire_config  (autofire_config),
      .cd32pad          (cd32pad),
      .usrrst           (usrrst),
      .cpurst           (cpurst),
      .cpuhlt           (cpuhlt),
      .fifo_full        (fifo_full),
      .host_cs          (host_cs),
      .host_adr         (host_adr),
      .host_we          (host_we),
      .host_bs          (host_bs),
      .host_wdat        (host_wdat),
      .host_rdat        (host_rdat),
      .host_ack         (host_ack)
      );

endmodule
